`timescale 1ns/1ps

module alu_test;


reg[31:0] instruction, regA, regB; 
// the address of regA is 00000, the address of regB is 00001
wire[31:0] result;
wire[2:0] flags; 
reg[39:0] name;

alu testalu(instruction, regA, regB, result, flags);

initial
begin

$display("instruction | name | regA | regB | result | flags");
$monitor("%b | %s | %b | %b | %b | %b",
instruction, name, regA, regB, result, flags);



#10 //add: flags[2] = 1'b1
instruction <= 32'b000000_00000_00001_00000_00000_100000;
regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
regB <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
name <= "add";

#10 //addu: result = 32'b0111_1111_1111_1111_1111_1111_1111_1111
instruction <= 32'b000000_00000_00001_00000_00000_100001;
regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
regB <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
name <= "addu";

#10 //addi: flags[2] = 1'b1
instruction <= 32'b001000_00001_00000_0000000000000001;
regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
regB <= 32'b0111_1111_1111_1111_1111_1111_1111_1111;
name <= "addi";

#10 //addiu: result = 32'b1000_0000_0000_0000_0000_0000_0000_0000
instruction <= 32'b001001_00001_00000_0000000000000001;
regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
regB <= 32'b0111_1111_1111_1111_1111_1111_1111_1111;
name <= "addiu";

#10 //sub: flags[2] = 1'b0
instruction <= 32'b000000_00000_00001_00000_00000_100010;
regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
regB <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
name <= "sub";

#10 //subu: result = 32'b0111_1111_1111_1111_1111_1111_1111_1111;
instruction <= 32'b000000_00000_00001_00000_00000_100011;
regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
regB <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
name <= "subu";

#10 //and: result = 32'b0000_0000_1111_0000_0000_0000_0000_1111;
instruction <= 32'b000000_00000_00001_00000_00000_100100;
regA <= 32'b0000_1111_1111_0000_0000_1111_1111_1111;
regB <= 32'b1111_0000_1111_1111_0000_0000_0000_1111;
name <= "and";

#10 //andi: result = 32'b0000_0000_0000_0000_1111_1111_1111_1111;
instruction <= 32'b001100_00000_00001_1111111111111111;
regA <= 32'b1111_1111_1111_1111_1111_1111_1111_1111;
regB <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
name <= "andi";

#10 //nor: result = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
instruction <= 32'b000000_00000_00001_00000_00000_100111;
regA <= 32'b1111_1111_1111_0000_0000_1111_1111_1111;
regB <= 32'b0000_0000_0000_0000_0000_1111_1111_1111;
name <= "nor";

#10 //or: result = 32'b1111_1111_1111_0000_0000_1111_1111_1111;
instruction <= 32'b000000_00000_00001_00000_00000_100101;
regA <= 32'b1111_1111_1111_0000_0000_1111_1111_1111;
regB <= 32'b0000_0000_0000_0000_0000_1111_1111_1111;

#10 //ori: result = 32'b0000_0000_0000_0000_1111_1111_1111_1111;
instruction <= 32'b001101_00000_00001_1111111111111111;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
regB <= 32'b0000_0000_0000_0000_0000_1111_1111_1111;
name <= "ori";

#10 //xor: result = 32'b1111_1111_1111_0000_0000_0000_0000_0000;
instruction <= 32'b000000_00000_00001_00000_00000_100110;
regA <= 32'b1111_1111_1111_0000_0000_1111_1111_1111;
regB <= 32'b0000_0000_0000_0000_0000_1111_1111_1111;
name <= "xor";

#10 //xori: result = 32'b1111_1111_1111_0000_0000_1111_1111_0000;
instruction <= 32'b001110_00000_00001_0000000000001111;
regA <= 32'b1111_1111_1111_0000_0000_1111_1111_1111;
regB <= 32'b0000_0000_0000_0000_0000_1111_1111_1111;
name <= "xori";

#10 //beq: tags[0] = 1'b1;
instruction <= 32'b000100_00000_00001_0000000000001111;
regA <= 32'b1111_1111_1111_0000_0000_1111_1111_1111;
regB <= 32'b1111_1111_1111_0000_0000_1111_1111_1111;
name <= "beq";

#10 //bne: tags[0] = 1'b1;
instruction <= 32'b000101_00000_00001_0000000000001111;
regA <= 32'b1111_1111_1111_0000_0000_1111_1111_1111;
regB <= 32'b1111_1111_1111_0000_0000_1111_1111_1110;
name <= "bne";

#10 //slt: tags[1] = 1'b1;
instruction <= 32'b000000_00000_00001_00000_00000_101010;
regA <= 32'b1111_1111_1111_0000_0000_1111_1111_1110;
regB <= 32'b1111_1111_1111_0000_0000_1111_1111_1111;
name <= "slt";

#10 //sltu: tags[1] = 1'b1;
instruction <= 32'b000000_00000_00001_00000_00000_101011;
regA <= 32'b1111_1111_1111_0000_0000_1111_1111_1110;
regB <= 32'b1111_1111_1111_0000_0000_1111_1111_1111;
name <= "sltu";

#10 //slti: tags[1] = 1'b0;
instruction <= 32'b001010_00000_00001_1000000000101011;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_1111;
regB <= 32'b1000_0000_0000_0000_0000_0000_0000_1111;
name <= "slti";

#10 //sltiu: tags[1] = 1'b1;
instruction <= 32'b001011_00000_00001_0000000000101011;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_1111;
regB <= 32'b1000_0000_0000_0000_0000_0000_0000_1111;
name <= "sltiu";

#10 //lw: result = 32'b0000_0000_0000_0000_0000_0000_0000_1111
instruction <= 32'b100011_00000_00001_0000000000000000;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_1111;
regB <= 32'b1000_0000_0000_0000_0000_0000_0000_1111;
name <= "lw";

#10 //sw: result = 32'b1000_0000_0000_0000_0000_0000_0000_1111
instruction <= 32'b101011_00001_00000_0000000000000000;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_1111;
regB <= 32'b1000_0000_0000_0000_0000_0000_0000_1111;
name <= "sw";

#10 //sll: result = 32'b1111_1111_0000_0000_1111_1111_1111_0000
instruction <= 32'b000000_00000_00001_00000_00100_000000;
regA <= 32'b1111_1111_1111_0000_0000_1111_1111_1110;
regB <= 32'b1111_1111_1111_0000_0000_1111_1111_1111;
name <= "sll";

#10 //sllv: result = 32'b1111_0000_0000_1111_1111_1111_0000_0000
instruction <= 32'b000000_00000_00001_00000_00100_000100;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_1000;
regB <= 32'b1111_1111_1111_0000_0000_1111_1111_1111;
name <= "sllv";

#10 //sra: result = 32'b1111_1111_1111_1111_0000_0000_1111_1111
instruction <= 32'b000000_00000_00001_00000_00100_000011;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_1000;
regB <= 32'b1111_1111_1111_0000_0000_1111_1111_1111;
name <= "sra";

#10 //srav: result = 32'b1111_1111_1111_1111_1111_0000_0000_1111
instruction <= 32'b000000_00000_00001_00000_00100_000111;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_1000;
regB <= 32'b1111_1111_1111_0000_0000_1111_1111_1111;
name <= "srav";

#10 //srl: result = 32'b0000_1111_1111_1111_0000_0000_1111_1111
instruction <= 32'b000000_00000_00001_00000_00100_000010;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_1000;
regB <= 32'b1111_1111_1111_0000_0000_1111_1111_1111;
name <= "srl";

#10 //srlv: result = 32'b0000_0000_1111_1111_1111_0000_0000_1111
instruction <= 32'b000000_00000_00001_00000_00100_000110;
regA <= 32'b0000_0000_0000_0000_0000_0000_0000_1000;
regB <= 32'b1111_1111_1111_0000_0000_1111_1111_1111;
name <= "srlv";

#10 $finish;
end

/*iverilog */
initial
begin            
    $dumpfile("wave.vcd");        
    $dumpvars(0, alu_test);    
end
/*iverilog */

endmodule